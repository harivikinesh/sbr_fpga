// fpu.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module fpu (
		input  wire [31:0] dataa,  // s1.dataa
		input  wire [31:0] datab,  //   .datab
		input  wire [3:0]  n,      //   .n
		output wire [31:0] result  //   .result
	);

	fpoint2_combi #(
		.arithmetic_present (1),
		.comparison_present (1)
	) nios_custom_instr_floating_point_2_combi_0 (
		.dataa  (dataa),  // s1.dataa
		.datab  (datab),  //   .datab
		.n      (n),      //   .n
		.result (result)  //   .result
	);

endmodule
